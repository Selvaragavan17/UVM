class seq_item extends uvm_sequence_item;
  rand bit [3:0]a;
  rand bit [3:0]b;
  rand bit [2:0]sel;
  rand bit [5:0]result;
  
  `uvm_objects_utils(seq_item);
  
  function new (string name="seq_item");
    super.new(name);
  endfunction
  
endclass
