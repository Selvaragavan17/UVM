interface intf(intput clk);
  logic clk;
  logic [3:0]a,b;
  logic [2:0]sel;
  logic [5:0]result;
endinterface
